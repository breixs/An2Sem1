library verilog;
use verilog.vl_types.all;
entity TransformNumber_tb is
end TransformNumber_tb;
