library verilog;
use verilog.vl_types.all;
entity transform_tb is
end transform_tb;
