module comp(input[7:0] in_0, input[7:0] in_1, output reg eq, output reg[7:0] max); reg [7:0] aux; initial begin eq=0; max=8'b10110100; end always@(in_1) begin aux=in_1; if (aux[7]==1) begin aux[7]=0; aux=~aux; aux=aux+1; end if(aux>in_0) begin max=aux; end else begin max=in_0; if(aux==in_0) begin max=8'b100000001; end end endmodule module comp_tb; reg[7:0] in_0; reg[7:0] in_1; wire eq; wire[7:0] max; comp uut(.in_0(in_0), .in_1(in_1), .eq(eq), .max(max)); integer k; initial begin $monitor("in_0=%8b, in_1=%8b\t\teq=%1b\tmax=%8b", in_0, in_1, eq, max); for(k = 0; k < 65536; k = k + 1) begin {in_0, in_1} = k; #1; end end endmodule
