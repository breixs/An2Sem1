library verilog;
use verilog.vl_types.all;
entity comp_tb is
end comp_tb;
