library verilog;
use verilog.vl_types.all;
entity nuj_tb is
end nuj_tb;
