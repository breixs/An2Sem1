library verilog;
use verilog.vl_types.all;
entity order_tb is
end order_tb;
