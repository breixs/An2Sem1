library verilog;
use verilog.vl_types.all;
entity diagram_tb is
end diagram_tb;
