module exercitiu 2
